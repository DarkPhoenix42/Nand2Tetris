LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY inc32_tb IS
END ENTITY;

ARCHITECTURE testbench OF inc32_tb IS
    COMPONENT inc32
        PORT (
            a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            o : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
        );
    END COMPONENT;

    SIGNAL a : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL o : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
    uut : inc32
    PORT MAP(
        a => a,
        o => o
    );
    PROCESS
    BEGIN
        a <= "00000000000000000000000000000000";
        WAIT FOR 10 us;
        ASSERT o = "00000000000000000000000000000001" REPORT "Test 1 failed" SEVERITY error;

        a <= "11111111111111111111111111111111";
        WAIT FOR 10 us;
        ASSERT o = "00000000000000000000000000000000" REPORT "Test 2 failed" SEVERITY error;

        WAIT;
    END PROCESS;
END ARCHITECTURE;